-- M�nica Colomera
-- M�dulo RAM 
-- Vers�o 0.1
--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ram is
    Port ( clk : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           addr : in  STD_LOGIC_VECTOR (7 downto 0);
           din : in  STD_LOGIC_VECTOR (7 downto 0);
           rw : in  STD_LOGIC;
           dout : out  STD_LOGIC_VECTOR (7 downto 0));
end ram;

architecture Behavioral of ram is

begin


end Behavioral;

